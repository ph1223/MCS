*****Example for including .vec file as input pattern****** 
.TITLE Current_mode_SA
*****************************
**     Library setting     **
*****************************
.protect
.include "/RAID2/COURSE/mcs/mcs020/Technology_files/7nm_TT.pm"
.unprotect

***************************************
**           Input vector            **
***************************************
.VEC 'input.vec'

*****************************
**     Voltage Source      **
*****************************
.global VDD GND

Vvdd VDD GND 0.7v
VWL  WLL  GND 0v

*****************************
**   Circuit Description   **
*****************************
.subckt inverter vin vout
Mp  vout  vin  VDD  x  pmos_sram  m=1
Mn  vout  vin  GND  x  nmos_sram  m=1
.ends

.subckt SRAM WL BL BLB
Mpr	 q	 qb  VDD  x  pmos_sram  m=1
Mnr  q   qb  GND  x  nmos_sram  m=1

Mpl  qb  q  VDD  x  pmos_sram  m=1
Mnl  qb  q  GND  x  nmos_sram  m=1

Mnpr BL  WL  q    x  nmos_sram  m=1
Mnpl BLB WL  qb   x  nmos_sram  m=1
.ends

.subckt SA BL BLB SEN output outputb
Mp1   outputb  SEN 	   VDD  x  pmos_sram  m=1
Mp2   output   SEN     VDD  x  pmos_sram  m=1
Mp3   outputb  output  VDD  x  pmos_sram  m=1
Mp4   output   outputb VDD  x  pmos_sram  m=1
Mn1   outputb  output   n1  x  nmos_sram  m=1
Mn2   output   outputb  n2  x  nmos_sram  m=1    
Mn3       n1   BL       n3  x  nmos_sram  m=1
Mn4       n2   BLB      n3  x  nmos_sram  m=1
Mn5       n3   SEN     GND  x  nmos_sram  m=1
.ends

Mp5   BL   pre     VDD  x  pmos_sram  m=1
Mp6   BLB  pre     VDD  x  pmos_sram  m=1
Mp7   BLB  pre      BL  x  pmos_sram  m=1

X0  	WL0	BL	BLB	SRAM
X1  	WLL	BL	BLB	SRAM
X2  	WLL	BL	BLB	SRAM
X3  	WLL	BL	BLB	SRAM
X4  	WLL	BL	BLB	SRAM
X5  	WLL	BL	BLB	SRAM
X6  	WLL	BL	BLB	SRAM
X7  	WLL	BL	BLB	SRAM
X8  	WLL	BL	BLB	SRAM
X9  	WLL	BL	BLB	SRAM
X10  	WLL	BL	BLB	SRAM
X11  	WLL	BL	BLB	SRAM
X12  	WLL	BL	BLB	SRAM
X13  	WLL	BL	BLB	SRAM
X14  	WLL	BL	BLB	SRAM
X15  	WLL	BL	BLB	SRAM

X16  	WLL	BL	BLB	SRAM
X17  	WLL	BL	BLB	SRAM
X18  	WLL	BL	BLB	SRAM
X19  	WLL	BL	BLB	SRAM
X20  	WLL	BL	BLB	SRAM
X21  	WLL	BL	BLB	SRAM
X22  	WLL	BL	BLB	SRAM
X23  	WLL	BL	BLB	SRAM
X24  	WLL	BL	BLB	SRAM
X25  	WLL	BL	BLB	SRAM
X26  	WLL	BL	BLB	SRAM
X27  	WLL	BL	BLB	SRAM
X28  	WLL	BL	BLB	SRAM
X29  	WLL	BL	BLB	SRAM
X30  	WLL	BL	BLB	SRAM
X31  	WLL	BL	BLB	SRAM

X32  	WLL	BL	BLB	SRAM
X33  	WLL	BL	BLB	SRAM
X34  	WLL	BL	BLB	SRAM
X35  	WLL	BL	BLB	SRAM
X36  	WLL	BL	BLB	SRAM
X37  	WLL	BL	BLB	SRAM
X38  	WLL	BL	BLB	SRAM
X39  	WLL	BL	BLB	SRAM
X40  	WLL	BL	BLB	SRAM
X41  	WLL	BL	BLB	SRAM
X42  	WLL	BL	BLB	SRAM
X43  	WLL	BL	BLB	SRAM
X44  	WLL	BL	BLB	SRAM
X45  	WLL	BL	BLB	SRAM
X46  	WLL	BL	BLB	SRAM
X47  	WLL	BL	BLB	SRAM

X48  	WLL	BL	BLB	SRAM
X49  	WLL	BL	BLB	SRAM
X50  	WLL	BL	BLB	SRAM
X51  	WLL	BL	BLB	SRAM
X52  	WLL	BL	BLB	SRAM
X53  	WLL	BL	BLB	SRAM
X54  	WLL	BL	BLB	SRAM
X55  	WLL	BL	BLB	SRAM
X56  	WLL	BL	BLB	SRAM
X57  	WLL	BL	BLB	SRAM
X58  	WLL	BL	BLB	SRAM
X59  	WLL	BL	BLB	SRAM
X60  	WLL	BL	BLB	SRAM
X61  	WLL	BL	BLB	SRAM
X62  	WLL	BL	BLB	SRAM
X63  	WLL	BL	BLB	SRAM

X64  	WLL	BL	BLB	SRAM
X65  	WLL	BL	BLB	SRAM
X66  	WLL	BL	BLB	SRAM
X67  	WLL	BL	BLB	SRAM
X68  	WLL	BL	BLB	SRAM
X69  	WLL	BL	BLB	SRAM
X70  	WLL	BL	BLB	SRAM
X71  	WLL	BL	BLB	SRAM
X72  	WLL	BL	BLB	SRAM
X73  	WLL	BL	BLB	SRAM
X74  	WLL	BL	BLB	SRAM
X75  	WLL	BL	BLB	SRAM
X76  	WLL	BL	BLB	SRAM
X77  	WLL	BL	BLB	SRAM
X78  	WLL	BL	BLB	SRAM
X79  	WLL	BL	BLB	SRAM

X80  	WLL	BL	BLB	SRAM
X81  	WLL	BL	BLB	SRAM
X82  	WLL	BL	BLB	SRAM
X83  	WLL	BL	BLB	SRAM
X84  	WLL	BL	BLB	SRAM
X85  	WLL	BL	BLB	SRAM
X86  	WLL	BL	BLB	SRAM
X87  	WLL	BL	BLB	SRAM
X88  	WLL	BL	BLB	SRAM
X89  	WLL	BL	BLB	SRAM
X90  	WLL	BL	BLB	SRAM
X91  	WLL	BL	BLB	SRAM
X92  	WLL	BL	BLB	SRAM
X93  	WLL	BL	BLB	SRAM
X94  	WLL	BL	BLB	SRAM
X95  	WLL	BL	BLB	SRAM

X96  	WLL	BL	BLB	SRAM
X97  	WLL	BL	BLB	SRAM
X98  	WLL	BL	BLB	SRAM
X99  	WLL	BL	BLB	SRAM
X100  	WLL	BL	BLB	SRAM
X101  	WLL	BL	BLB	SRAM
X102  	WLL	BL	BLB	SRAM
X103  	WLL	BL	BLB	SRAM
X104  	WLL	BL	BLB	SRAM
X105  	WLL	BL	BLB	SRAM
X106  	WLL	BL	BLB	SRAM
X107  	WLL	BL	BLB	SRAM
X108  	WLL	BL	BLB	SRAM
X109  	WLL	BL	BLB	SRAM
X110  	WLL	BL	BLB	SRAM
X111  	WLL	BL	BLB	SRAM

X112  	WLL	BL	BLB	SRAM
X113  	WLL	BL	BLB	SRAM
X114  	WLL	BL	BLB	SRAM
X115  	WLL	BL	BLB	SRAM
X116  	WLL	BL	BLB	SRAM
X117  	WLL	BL	BLB	SRAM
X118  	WLL	BL	BLB	SRAM
X119  	WLL	BL	BLB	SRAM
X120  	WLL	BL	BLB	SRAM
X121  	WLL	BL	BLB	SRAM
X122  	WLL	BL	BLB	SRAM
X123  	WLL	BL	BLB	SRAM
X124  	WLL	BL	BLB	SRAM
X125  	WLL	BL	BLB	SRAM
X126  	WLL	BL	BLB	SRAM
X127  	WLL	BL	BLB	SRAM

X128  	WLL	BL	BLB	SRAM
X129  	WLL	BL	BLB	SRAM
X130  	WLL	BL	BLB	SRAM
X131  	WLL	BL	BLB	SRAM
X132  	WLL	BL	BLB	SRAM
X133  	WLL	BL	BLB	SRAM
X134  	WLL	BL	BLB	SRAM
X135  	WLL	BL	BLB	SRAM
X136  	WLL	BL	BLB	SRAM
X137  	WLL	BL	BLB	SRAM
X138  	WLL	BL	BLB	SRAM
X139  	WLL	BL	BLB	SRAM
X140  	WLL	BL	BLB	SRAM
X141  	WLL	BL	BLB	SRAM
X142  	WLL	BL	BLB	SRAM
X143  	WLL	BL	BLB	SRAM

X144  	WLL	BL	BLB	SRAM
X145  	WLL	BL	BLB	SRAM
X146  	WLL	BL	BLB	SRAM
X147  	WLL	BL	BLB	SRAM
X148  	WLL	BL	BLB	SRAM
X149  	WLL	BL	BLB	SRAM
X150  	WLL	BL	BLB	SRAM
X151  	WLL	BL	BLB	SRAM
X152  	WLL	BL	BLB	SRAM
X153  	WLL	BL	BLB	SRAM
X154  	WLL	BL	BLB	SRAM
X155  	WLL	BL	BLB	SRAM
X156  	WLL	BL	BLB	SRAM
X157  	WLL	BL	BLB	SRAM
X158  	WLL	BL	BLB	SRAM
X159  	WLL	BL	BLB	SRAM

X160  	WLL	BL	BLB	SRAM
X161  	WLL	BL	BLB	SRAM
X162  	WLL	BL	BLB	SRAM
X163  	WLL	BL	BLB	SRAM
X164  	WLL	BL	BLB	SRAM
X165  	WLL	BL	BLB	SRAM
X166  	WLL	BL	BLB	SRAM
X167  	WLL	BL	BLB	SRAM
X168  	WLL	BL	BLB	SRAM
X169  	WLL	BL	BLB	SRAM
X170  	WLL	BL	BLB	SRAM
X171  	WLL	BL	BLB	SRAM
X172  	WLL	BL	BLB	SRAM
X173  	WLL	BL	BLB	SRAM
X174  	WLL	BL	BLB	SRAM
X175  	WLL	BL	BLB	SRAM

X176  	WLL	BL	BLB	SRAM
X177  	WLL	BL	BLB	SRAM
X178  	WLL	BL	BLB	SRAM
X179  	WLL	BL	BLB	SRAM
X180  	WLL	BL	BLB	SRAM
X181  	WLL	BL	BLB	SRAM
X182  	WLL	BL	BLB	SRAM
X183  	WLL	BL	BLB	SRAM
X184  	WLL	BL	BLB	SRAM
X185  	WLL	BL	BLB	SRAM
X186  	WLL	BL	BLB	SRAM
X187  	WLL	BL	BLB	SRAM
X188  	WLL	BL	BLB	SRAM
X189  	WLL	BL	BLB	SRAM
X190  	WLL	BL	BLB	SRAM
X191  	WLL	BL	BLB	SRAM

X192  	WLL	BL	BLB	SRAM
X193  	WLL	BL	BLB	SRAM
X194  	WLL	BL	BLB	SRAM
X195  	WLL	BL	BLB	SRAM
X196  	WLL	BL	BLB	SRAM
X197  	WLL	BL	BLB	SRAM
X198  	WLL	BL	BLB	SRAM
X199  	WLL	BL	BLB	SRAM
X200  	WLL	BL	BLB	SRAM
X201  	WLL	BL	BLB	SRAM
X202  	WLL	BL	BLB	SRAM
X203  	WLL	BL	BLB	SRAM
X204  	WLL	BL	BLB	SRAM
X205  	WLL	BL	BLB	SRAM
X206  	WLL	BL	BLB	SRAM
X207  	WLL	BL	BLB	SRAM

X208  	WLL	BL	BLB	SRAM
X209  	WLL	BL	BLB	SRAM
X210  	WLL	BL	BLB	SRAM
X211  	WLL	BL	BLB	SRAM
X212  	WLL	BL	BLB	SRAM
X213  	WLL	BL	BLB	SRAM
X214  	WLL	BL	BLB	SRAM
X215  	WLL	BL	BLB	SRAM
X216  	WLL	BL	BLB	SRAM
X217  	WLL	BL	BLB	SRAM
X218  	WLL	BL	BLB	SRAM
X219  	WLL	BL	BLB	SRAM
X220  	WLL	BL	BLB	SRAM
X221  	WLL	BL	BLB	SRAM
X222  	WLL	BL	BLB	SRAM
X223  	WLL	BL	BLB	SRAM

X224  	WLL	BL	BLB	SRAM
X225  	WLL	BL	BLB	SRAM
X226  	WLL	BL	BLB	SRAM
X227  	WLL	BL	BLB	SRAM
X228  	WLL	BL	BLB	SRAM
X229  	WLL	BL	BLB	SRAM
X230  	WLL	BL	BLB	SRAM
X231  	WLL	BL	BLB	SRAM
X232  	WLL	BL	BLB	SRAM
X233  	WLL	BL	BLB	SRAM
X234  	WLL	BL	BLB	SRAM
X235  	WLL	BL	BLB	SRAM
X236  	WLL	BL	BLB	SRAM
X237  	WLL	BL	BLB	SRAM
X238  	WLL	BL	BLB	SRAM
X239  	WLL	BL	BLB	SRAM

X240  	WLL	BL	BLB	SRAM
X241  	WLL	BL	BLB	SRAM
X242  	WLL	BL	BLB	SRAM
X243  	WLL	BL	BLB	SRAM
X244  	WLL	BL	BLB	SRAM
X245  	WLL	BL	BLB	SRAM
X246  	WLL	BL	BLB	SRAM
X247  	WLL	BL	BLB	SRAM
X248  	WLL	BL	BLB	SRAM
X249  	WLL	BL	BLB	SRAM
X250  	WLL	BL	BLB	SRAM
X251  	WLL	BL	BLB	SRAM
X252  	WLL	BL	BLB	SRAM
X253  	WLL	BL	BLB	SRAM
X254  	WLL	BL	BLB	SRAM
X255  	WLL	BL	BLB	SRAM

X256  	WLL	BL	BLB	SRAM
X257  	WLL	BL	BLB	SRAM
X258  	WLL	BL	BLB	SRAM
X259  	WLL	BL	BLB	SRAM
X260  	WLL	BL	BLB	SRAM
X261  	WLL	BL	BLB	SRAM
X262  	WLL	BL	BLB	SRAM
X263  	WLL	BL	BLB	SRAM
X264  	WLL	BL	BLB	SRAM
X265  	WLL	BL	BLB	SRAM
X266  	WLL	BL	BLB	SRAM
X267  	WLL	BL	BLB	SRAM
X268  	WLL	BL	BLB	SRAM
X269  	WLL	BL	BLB	SRAM
X270  	WLL	BL	BLB	SRAM
X271  	WLL	BL	BLB	SRAM

X272  	WLL	BL	BLB	SRAM
X273  	WLL	BL	BLB	SRAM
X274  	WLL	BL	BLB	SRAM
X275  	WLL	BL	BLB	SRAM
X276  	WLL	BL	BLB	SRAM
X277  	WLL	BL	BLB	SRAM
X278  	WLL	BL	BLB	SRAM
X279  	WLL	BL	BLB	SRAM
X280  	WLL	BL	BLB	SRAM
X281  	WLL	BL	BLB	SRAM
X282  	WLL	BL	BLB	SRAM
X283  	WLL	BL	BLB	SRAM
X284  	WLL	BL	BLB	SRAM
X285  	WLL	BL	BLB	SRAM
X286  	WLL	BL	BLB	SRAM
X287  	WLL	BL	BLB	SRAM

X288  	WLL	BL	BLB	SRAM
X289  	WLL	BL	BLB	SRAM
X290  	WLL	BL	BLB	SRAM
X291  	WLL	BL	BLB	SRAM
X292  	WLL	BL	BLB	SRAM
X293  	WLL	BL	BLB	SRAM
X294  	WLL	BL	BLB	SRAM
X295  	WLL	BL	BLB	SRAM
X296  	WLL	BL	BLB	SRAM
X297  	WLL	BL	BLB	SRAM
X298  	WLL	BL	BLB	SRAM
X299  	WLL	BL	BLB	SRAM
X300  	WLL	BL	BLB	SRAM
X301  	WLL	BL	BLB	SRAM
X302  	WLL	BL	BLB	SRAM
X303  	WLL	BL	BLB	SRAM

X304  	WLL	BL	BLB	SRAM
X305  	WLL	BL	BLB	SRAM
X306  	WLL	BL	BLB	SRAM
X307  	WLL	BL	BLB	SRAM
X308  	WLL	BL	BLB	SRAM
X309  	WLL	BL	BLB	SRAM
X310  	WLL	BL	BLB	SRAM
X311  	WLL	BL	BLB	SRAM
X312  	WLL	BL	BLB	SRAM
X313  	WLL	BL	BLB	SRAM
X314  	WLL	BL	BLB	SRAM
X315  	WLL	BL	BLB	SRAM
X316  	WLL	BL	BLB	SRAM
X317  	WLL	BL	BLB	SRAM
X318  	WLL	BL	BLB	SRAM
X319  	WLL	BL	BLB	SRAM

X320  	WLL	BL	BLB	SRAM
X321  	WLL	BL	BLB	SRAM
X322  	WLL	BL	BLB	SRAM
X323  	WLL	BL	BLB	SRAM
X324  	WLL	BL	BLB	SRAM
X325  	WLL	BL	BLB	SRAM
X326  	WLL	BL	BLB	SRAM
X327  	WLL	BL	BLB	SRAM
X328  	WLL	BL	BLB	SRAM
X329  	WLL	BL	BLB	SRAM
X330  	WLL	BL	BLB	SRAM
X331  	WLL	BL	BLB	SRAM
X332  	WLL	BL	BLB	SRAM
X333  	WLL	BL	BLB	SRAM
X334  	WLL	BL	BLB	SRAM
X335  	WLL	BL	BLB	SRAM

X336  	WLL	BL	BLB	SRAM
X337  	WLL	BL	BLB	SRAM
X338  	WLL	BL	BLB	SRAM
X339  	WLL	BL	BLB	SRAM
X340  	WLL	BL	BLB	SRAM
X341  	WLL	BL	BLB	SRAM
X342  	WLL	BL	BLB	SRAM
X343  	WLL	BL	BLB	SRAM
X344  	WLL	BL	BLB	SRAM
X345  	WLL	BL	BLB	SRAM
X346  	WLL	BL	BLB	SRAM
X347  	WLL	BL	BLB	SRAM
X348  	WLL	BL	BLB	SRAM
X349  	WLL	BL	BLB	SRAM
X350  	WLL	BL	BLB	SRAM
X351  	WLL	BL	BLB	SRAM

X352  	WLL	BL	BLB	SRAM
X353  	WLL	BL	BLB	SRAM
X354  	WLL	BL	BLB	SRAM
X355  	WLL	BL	BLB	SRAM
X356  	WLL	BL	BLB	SRAM
X357  	WLL	BL	BLB	SRAM
X358  	WLL	BL	BLB	SRAM
X359  	WLL	BL	BLB	SRAM
X360  	WLL	BL	BLB	SRAM
X361  	WLL	BL	BLB	SRAM
X362  	WLL	BL	BLB	SRAM
X363  	WLL	BL	BLB	SRAM
X364  	WLL	BL	BLB	SRAM
X365  	WLL	BL	BLB	SRAM
X366  	WLL	BL	BLB	SRAM
X367  	WLL	BL	BLB	SRAM

X368  	WLL	BL	BLB	SRAM
X369  	WLL	BL	BLB	SRAM
X370  	WLL	BL	BLB	SRAM
X371  	WLL	BL	BLB	SRAM
X372  	WLL	BL	BLB	SRAM
X373  	WLL	BL	BLB	SRAM
X374  	WLL	BL	BLB	SRAM
X375  	WLL	BL	BLB	SRAM
X376  	WLL	BL	BLB	SRAM
X377  	WLL	BL	BLB	SRAM
X378  	WLL	BL	BLB	SRAM
X379  	WLL	BL	BLB	SRAM
X380  	WLL	BL	BLB	SRAM
X381  	WLL	BL	BLB	SRAM
X382  	WLL	BL	BLB	SRAM
X383  	WLL	BL	BLB	SRAM

X384  	WLL	BL	BLB	SRAM
X385  	WLL	BL	BLB	SRAM
X386  	WLL	BL	BLB	SRAM
X387  	WLL	BL	BLB	SRAM
X388  	WLL	BL	BLB	SRAM
X389  	WLL	BL	BLB	SRAM
X390  	WLL	BL	BLB	SRAM
X391  	WLL	BL	BLB	SRAM
X392  	WLL	BL	BLB	SRAM
X393  	WLL	BL	BLB	SRAM
X394  	WLL	BL	BLB	SRAM
X395  	WLL	BL	BLB	SRAM
X396  	WLL	BL	BLB	SRAM
X397  	WLL	BL	BLB	SRAM
X398  	WLL	BL	BLB	SRAM
X399  	WLL	BL	BLB	SRAM

X400  	WLL	BL	BLB	SRAM
X401  	WLL	BL	BLB	SRAM
X402  	WLL	BL	BLB	SRAM
X403  	WLL	BL	BLB	SRAM
X404  	WLL	BL	BLB	SRAM
X405  	WLL	BL	BLB	SRAM
X406  	WLL	BL	BLB	SRAM
X407  	WLL	BL	BLB	SRAM
X408  	WLL	BL	BLB	SRAM
X409  	WLL	BL	BLB	SRAM
X410  	WLL	BL	BLB	SRAM
X411  	WLL	BL	BLB	SRAM
X412  	WLL	BL	BLB	SRAM
X413  	WLL	BL	BLB	SRAM
X414  	WLL	BL	BLB	SRAM
X415  	WLL	BL	BLB	SRAM

X416  	WLL	BL	BLB	SRAM
X417  	WLL	BL	BLB	SRAM
X418  	WLL	BL	BLB	SRAM
X419  	WLL	BL	BLB	SRAM
X420  	WLL	BL	BLB	SRAM
X421  	WLL	BL	BLB	SRAM
X422  	WLL	BL	BLB	SRAM
X423  	WLL	BL	BLB	SRAM
X424  	WLL	BL	BLB	SRAM
X425  	WLL	BL	BLB	SRAM
X426  	WLL	BL	BLB	SRAM
X427  	WLL	BL	BLB	SRAM
X428  	WLL	BL	BLB	SRAM
X429  	WLL	BL	BLB	SRAM
X430  	WLL	BL	BLB	SRAM
X431  	WLL	BL	BLB	SRAM

X432  	WLL	BL	BLB	SRAM
X433  	WLL	BL	BLB	SRAM
X434  	WLL	BL	BLB	SRAM
X435  	WLL	BL	BLB	SRAM
X436  	WLL	BL	BLB	SRAM
X437  	WLL	BL	BLB	SRAM
X438  	WLL	BL	BLB	SRAM
X439  	WLL	BL	BLB	SRAM
X440  	WLL	BL	BLB	SRAM
X441  	WLL	BL	BLB	SRAM
X442  	WLL	BL	BLB	SRAM
X443  	WLL	BL	BLB	SRAM
X444  	WLL	BL	BLB	SRAM
X445  	WLL	BL	BLB	SRAM
X446  	WLL	BL	BLB	SRAM
X447  	WLL	BL	BLB	SRAM

X448  	WLL	BL	BLB	SRAM
X449  	WLL	BL	BLB	SRAM
X450  	WLL	BL	BLB	SRAM
X451  	WLL	BL	BLB	SRAM
X452  	WLL	BL	BLB	SRAM
X453  	WLL	BL	BLB	SRAM
X454  	WLL	BL	BLB	SRAM
X455  	WLL	BL	BLB	SRAM
X456  	WLL	BL	BLB	SRAM
X457  	WLL	BL	BLB	SRAM
X458  	WLL	BL	BLB	SRAM
X459  	WLL	BL	BLB	SRAM
X460  	WLL	BL	BLB	SRAM
X461  	WLL	BL	BLB	SRAM
X462  	WLL	BL	BLB	SRAM
X463  	WLL	BL	BLB	SRAM

X464  	WLL	BL	BLB	SRAM
X465  	WLL	BL	BLB	SRAM
X466  	WLL	BL	BLB	SRAM
X467  	WLL	BL	BLB	SRAM
X468  	WLL	BL	BLB	SRAM
X469  	WLL	BL	BLB	SRAM
X470  	WLL	BL	BLB	SRAM
X471  	WLL	BL	BLB	SRAM
X472  	WLL	BL	BLB	SRAM
X473  	WLL	BL	BLB	SRAM
X474  	WLL	BL	BLB	SRAM
X475  	WLL	BL	BLB	SRAM
X476  	WLL	BL	BLB	SRAM
X477  	WLL	BL	BLB	SRAM
X478  	WLL	BL	BLB	SRAM
X479  	WLL	BL	BLB	SRAM

X480  	WLL	BL	BLB	SRAM
X481  	WLL	BL	BLB	SRAM
X482  	WLL	BL	BLB	SRAM
X483  	WLL	BL	BLB	SRAM
X484  	WLL	BL	BLB	SRAM
X485  	WLL	BL	BLB	SRAM
X486  	WLL	BL	BLB	SRAM
X487  	WLL	BL	BLB	SRAM
X488  	WLL	BL	BLB	SRAM
X489  	WLL	BL	BLB	SRAM
X490  	WLL	BL	BLB	SRAM
X491  	WLL	BL	BLB	SRAM
X492  	WLL	BL	BLB	SRAM
X493  	WLL	BL	BLB	SRAM
X494  	WLL	BL	BLB	SRAM
X495  	WLL	BL	BLB	SRAM

X496  	WLL	BL	BLB	SRAM
X497  	WLL	BL	BLB	SRAM
X498  	WLL	BL	BLB	SRAM
X499  	WLL	BL	BLB	SRAM
X500  	WLL	BL	BLB	SRAM
X501  	WLL	BL	BLB	SRAM
X502  	WLL	BL	BLB	SRAM
X503  	WLL	BL	BLB	SRAM
X504  	WLL	BL	BLB	SRAM
X505  	WLL	BL	BLB	SRAM
X506  	WLL	BL	BLB	SRAM
X507  	WLL	BL	BLB	SRAM
X508  	WLL	BL	BLB	SRAM
X509  	WLL	BL	BLB	SRAM
X510  	WLL	BL	BLB	SRAM
X511  	WLL	BL	BLB	SRAM

X512    BL  BLB SEN dout  doutb SA

*** wire loading/um
***	0.16fF/um     0.16*sqrt(0.027(um^2))=0.0263fF
***0.0263*512= 13.46fF
CBLB BLB GND 13.46fF
CBL   BL GND 13.46fF

.IC V(x0.q) = 0.7v

.op
.option post     
.options probe   
.probe v(*) i(*) 
.option captab   
.tran 0.01ns 10ns

.measure sensingtime
+ TRIG v(SEN) VAL='0.35' RISE=5
+ TARG v(doutb) VAL='0.01' FALL=5

.measure TRAN pwr avg power from=1n to=9n
.TEMP 25

.end